/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
creaded: 2017/6/6 
madified:
***********************************************/
// `include "axil_macro.sv"

// axi_stream_inf #(.DSIZE(8))  tx_udp_inf                         (.aclk(mac_clk_125M),.aresetn(mac_rst_n),.aclken(1'b1));
//
// `define DEF_COPY_AXIS(up_stream,name)\
