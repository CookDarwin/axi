/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2020-01-14 13:52:15 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module data_intc_M2S_force_robin#(
    parameter  NUM = 8
)(
    data_inf_c.slaver s00 [NUM-1:0],
    data_inf_c.master m00
);

//==========================================================================
//-------- define ----------------------------------------------------------
logic [$clog2(NUM)-1:0]  robin_index ;
logic from_up_vld;
logic to_up_ready;
//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
